module random_generator(
    output reg [0:
    );
    initial begin
    a = $urandom_rang(0, 10)

        case (a)

        endcase
    end
endmodule
