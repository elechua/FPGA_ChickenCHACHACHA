module next_turn(
    input clk, 
    input [2-1:0] N,
    input [2-1:0] T,
    input statecombo_next_turn,
    output [2-1:0] result
    // Q가 100에서 101
    // Q가 101에서 110으로 바뀌는 때가
    );
endmodule
