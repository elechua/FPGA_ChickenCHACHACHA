module random_generator(
    output reg random_order
);
    // 각 타일 위치를 몇비트로 설정하지 -> 6 bit => 24*6=144 bit?
    reg [23:0] orders [0:9]  // 일단은 10개만 
    reg [4:0] random_number;  // random number (0-9)
    
    initial begin
        orders[0] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[1] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[2] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[3] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[4] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[5] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[6] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[7] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[8] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
        orders[9] = 144'b000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000_000000;
    end // 첫번째 6bit 첫번째 그림 위치. 두번째 6비트 두번째 그림 위치 등으로 하면 될거같은데

    random_number <= $urandom % 10;  // random number (0-9)

    random_order <= order[random_number];

endmodule

