module control_unit(
    input clk, win, go, c,
    output Q, R, A, B
    );
    
endmodule
