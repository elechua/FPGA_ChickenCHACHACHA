module top_module(

    );
    
    control_unit cu(); //
    data_path dp(); //
    data_memory dm(); //
    random_generator rg(); // ��
endmodule
