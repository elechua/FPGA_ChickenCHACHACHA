module random_generator(
    input rst,
    output reg [96-1:0] random_edge_order
    output reg [48-1:0] random_center_order
);
    reg [96-1:0] edge_orders [0:9]  // 일단은 10개만 
    reg [48-1:0] center_orders [0:9]
    reg [4:0] random_number;  // random number (0-9)
    
    initial begin
        edge_orders[0] = 96'b1010_0001_0100_0011_0111_1001_0011_0010_0101_0111_0110_1011_0000_0001_1010_0100_0110_1000_1001_1011_1000_0000_0101_0010;
        edge_orders[1] = 96'b0001_0100_1010_0010_0011_1000_0111_0110_0101_1001_1000_0001_0000_1011_0000_0010_0011_0101_0111_1001_0100_1011_1010_0110;
        edge_orders[2] = 96'b0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011_0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011;
        edge_orders[3] = 96'b0001_1010_0010_0110_1000_0011_1011_0100_0001_0000_0110_1000_0011_1011_0111_1010_1001_0100_0000_0101_0010_0111_1001_0101;
        edge_orders[4] = 96'b1011_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1011_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000;
        edge_orders[5] = 96'b0000_0111_0001_0100_0011_1001_1010_0010_0110_0101_1000_1011_0000_0100_0011_0001_0111_0010_1001_1010_1011_0110_1000_0101;
        edge_orders[6] = 96'b0001_0110_0111_0010_0000_0100_0101_0110_0011_1010_1011_1001_0000_1010_0100_1000_0001_0111_1001_0011_0010_1011_1000_0101;
        edge_orders[7] = 96'b0010_1010_0111_1000_0101_0001_0100_1010_1001_0110_0000_0111_1011_0001_0000_0010_0110_1000_1001_0011_0100_1011_0101_0011;
        edge_orders[8] = 96'b0011_0110_0010_0100_0101_0001_0111_1000_0000_1001_1011_1010_0000_0100_0110_1011_0010_0011_0101_0111_1000_1010_0001_1001;
        edge_orders[9] = 96'b0110_1011_0000_0011_0010_0101_1001_0100_0001_1010_1000_1011_1001_0110_0011_0111_0000_1010_0010_1000_0101_0111_0100_0001;
        
        center_orders[0] = 48'b0000_0001_0010_0011_0100_0101_0110_0111_1000_1001_1010_1011;
        center_orders[1] = 48'b1011_1010_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000;
        center_orders[2] = 48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        center_orders[3] = 48'b0001_0111_0100_0000_1011_0101_0010_1000_1010_1001_0011_0110;
        center_orders[4] = 48'b0010_0001_1011_0000_0011_1010_0100_0101_1000_0111_1001_0110;
        center_orders[5] = 48'b0111_0000_0001_1000_0110_0101_1011_0100_1001_0010_1010_0011;
        center_orders[6] = 48'b1001_1000_0111_0001_0010_0000_0110_0011_1011_1010_0100_0101;
        center_orders[7] = 48'b0101_0000_0100_0110_0001_1011_1000_0111_0010_1001_0011_1010;
        center_orders[8] = 48'b0000_0010_0011_1011_0111_0001_1000_0110_1001_0100_1010_0101;
        center_orders[9] = 48'b0010_0111_0011_0110_0000_0101_0001_1000_1011_0100_1010_1001;

    end

    always @ (posedge rst) begin
        if (rst)
            random_number <= $urandom % 10;
    end

    //assign random_edge_order <= edge_order[random_number];
    //assign random_center_order <= center_order[random_number];

    assign random_edge_order <= edge_order[0];
    assign random_center_order <= center_order[0];
    
endmodule
